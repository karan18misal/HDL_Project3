module multiplier(input [15:0]a, input [15:0]b, output [31:0]y);
wire [31:0]y0;
wire [31:0]y1;
wire [31:0]y2;
wire [31:0]y3;
wire [31:0]y4;
wire [31:0]y5;
wire [31:0]y6;
wire [31:0]y7;
wire [31:0]y8;
wire [31:0]y9;
wire [31:0]y10;
wire [31:0]y11;
wire [31:0]y12;
wire [31:0]y13;
wire [31:0]y14;
wire [31:0]y15;

wire [31:0]s0;
wire [31:0]s1;
wire [31:0]s2;
wire [31:0]s3;
wire [31:0]s4;
wire [31:0]s5;
wire [31:0]s6;
wire [31:0]s7;
wire [31:0]s8;
wire [31:0]s9;
wire [31:0]s10;
wire [31:0]s11;
wire [31:0]s12;
wire [31:0]s13;
wire [31:0]s14;

wire cout0, cout1, cout2, cout3, cout4, cout5, cout6, cout7, cout8, cout9, cout10, cout11, cout12, cout13, cout14;

assign y0[0]  = a[0]  & b[0];
assign y0[1]  = a[1]  & b[0];
assign y0[2]  = a[2]  & b[0];
assign y0[3]  = a[3]  & b[0];
assign y0[4]  = a[4]  & b[0];
assign y0[5]  = a[5]  & b[0];
assign y0[6]  = a[6]  & b[0];
assign y0[7]  = a[7]  & b[0];
assign y0[8]  = a[8]  & b[0];
assign y0[9]  = a[9]  & b[0];
assign y0[10] = a[10] & b[0];
assign y0[11] = a[11] & b[0];
assign y0[12] = a[12] & b[0];
assign y0[13] = a[13] & b[0];
assign y0[14] = a[14] & b[0];
assign y0[15] = a[15] & b[0];
assign y0[31:16] = 16'b0;
  
assign y1[0]  = 1'b0;           
assign y1[1]  = a[0]  & b[1];
assign y1[2]  = a[1]  & b[1];
assign y1[3]  = a[2]  & b[1];
assign y1[4]  = a[3]  & b[1];
assign y1[5]  = a[4]  & b[1];
assign y1[6]  = a[5]  & b[1];
assign y1[7]  = a[6]  & b[1];
assign y1[8]  = a[7]  & b[1];
assign y1[9]  = a[8]  & b[1];
assign y1[10] = a[9]  & b[1];
assign y1[11] = a[10] & b[1];
assign y1[12] = a[11] & b[1];
assign y1[13] = a[12] & b[1];
assign y1[14] = a[13] & b[1];
assign y1[15] = a[14] & b[1];
assign y1[16] = a[15] & b[1];
assign y1[31:17] = 15'b0;
  
assign y2[1:0] = 2'b00;
assign y2[2]  = a[0]  & b[2];
assign y2[3]  = a[1]  & b[2];
assign y2[4]  = a[2]  & b[2];
assign y2[5]  = a[3]  & b[2];
assign y2[6]  = a[4]  & b[2];
assign y2[7]  = a[5]  & b[2];
assign y2[8]  = a[6]  & b[2];
assign y2[9]  = a[7]  & b[2];
assign y2[10] = a[8]  & b[2];
assign y2[11] = a[9]  & b[2];
assign y2[12] = a[10] & b[2];
assign y2[13] = a[11] & b[2];
assign y2[14] = a[12] & b[2];
assign y2[15] = a[13] & b[2];
assign y2[16] = a[14] & b[2];
assign y2[17] = a[15] & b[2];
assign y2[31:18] = 14'b0;
  
assign y3[2:0] = 3'b000;
assign y3[3]  = a[0]  & b[3];
assign y3[4]  = a[1]  & b[3];
assign y3[5]  = a[2]  & b[3];
assign y3[6]  = a[3]  & b[3];
assign y3[7]  = a[4]  & b[3];
assign y3[8]  = a[5]  & b[3];
assign y3[9]  = a[6]  & b[3];
assign y3[10] = a[7]  & b[3];
assign y3[11] = a[8]  & b[3];
assign y3[12] = a[9]  & b[3];
assign y3[13] = a[10] & b[3];
assign y3[14] = a[11] & b[3];
assign y3[15] = a[12] & b[3];
assign y3[16] = a[13] & b[3];
assign y3[17] = a[14] & b[3];
assign y3[18] = a[15] & b[3];
assign y3[31:19] = 13'b0;
  
assign y4[3:0] = 4'b0000;
assign y4[4]  = a[0]  & b[4];
assign y4[5]  = a[1]  & b[4];
assign y4[6]  = a[2]  & b[4];
assign y4[7]  = a[3]  & b[4];
assign y4[8]  = a[4]  & b[4];
assign y4[9]  = a[5]  & b[4];
assign y4[10] = a[6]  & b[4];
assign y4[11] = a[7]  & b[4];
assign y4[12] = a[8]  & b[4];
assign y4[13] = a[9]  & b[4];
assign y4[14] = a[10] & b[4];
assign y4[15] = a[11] & b[4];
assign y4[16] = a[12] & b[4];
assign y4[17] = a[13] & b[4];
assign y4[18] = a[14] & b[4];
assign y4[19] = a[15] & b[4];
assign y4[31:20] = 12'b0;

assign y5[4:0] = 5'b00000;
assign y5[5]  = a[0]  & b[5];
assign y5[6]  = a[1]  & b[5];
assign y5[7]  = a[2]  & b[5];
assign y5[8]  = a[3]  & b[5];
assign y5[9]  = a[4]  & b[5];
assign y5[10] = a[5]  & b[5];
assign y5[11] = a[6]  & b[5];
assign y5[12] = a[7]  & b[5];
assign y5[13] = a[8]  & b[5];
assign y5[14] = a[9]  & b[5];
assign y5[15] = a[10] & b[5];
assign y5[16] = a[11] & b[5];
assign y5[17] = a[12] & b[5];
assign y5[18] = a[13] & b[5];
assign y5[19] = a[14] & b[5];
assign y5[20] = a[15] & b[5];
assign y5[31:21] = 11'b0;

assign y6[5:0] = 6'b0;
assign y6[6]  = a[0]  & b[6];
assign y6[7]  = a[1]  & b[6];
assign y6[8]  = a[2]  & b[6];
assign y6[9]  = a[3]  & b[6];
assign y6[10] = a[4]  & b[6];
assign y6[11] = a[5]  & b[6];
assign y6[12] = a[6]  & b[6];
assign y6[13] = a[7]  & b[6];
assign y6[14] = a[8]  & b[6];
assign y6[15] = a[9]  & b[6];
assign y6[16] = a[10] & b[6];
assign y6[17] = a[11] & b[6];
assign y6[18] = a[12] & b[6];
assign y6[19] = a[13] & b[6];
assign y6[20] = a[14] & b[6];
assign y6[21] = a[15] & b[6];
assign y6[31:22] = 10'b0;

assign y7[6:0] = 7'b0;
assign y7[7]  = a[0]  & b[7];
assign y7[8]  = a[1]  & b[7];
assign y7[9]  = a[2]  & b[7];
assign y7[10] = a[3]  & b[7];
assign y7[11] = a[4]  & b[7];
assign y7[12] = a[5]  & b[7];
assign y7[13] = a[6]  & b[7];
assign y7[14] = a[7]  & b[7];
assign y7[15] = a[8]  & b[7];
assign y7[16] = a[9]  & b[7];
assign y7[17] = a[10] & b[7];
assign y7[18] = a[11] & b[7];
assign y7[19] = a[12] & b[7];
assign y7[20] = a[13] & b[7];
assign y7[21] = a[14] & b[7];
assign y7[22] = a[15] & b[7];
assign y7[31:23] = 9'b0;

assign y8[7:0] = 8'b0;
assign y8[8]  = a[0]  & b[8];
assign y8[9]  = a[1]  & b[8];
assign y8[10] = a[2]  & b[8];
assign y8[11] = a[3]  & b[8];
assign y8[12] = a[4]  & b[8];
assign y8[13] = a[5]  & b[8];
assign y8[14] = a[6]  & b[8];
assign y8[15] = a[7]  & b[8];
assign y8[16] = a[8]  & b[8];
assign y8[17] = a[9]  & b[8];
assign y8[18] = a[10] & b[8];
assign y8[19] = a[11] & b[8];
assign y8[20] = a[12] & b[8];
assign y8[21] = a[13] & b[8];
assign y8[22] = a[14] & b[8];
assign y8[23] = a[15] & b[8];
assign y8[31:24] = 8'b0;

assign y9[8:0] = 9'b0;
assign y9[9]  = a[0]  & b[9];
assign y9[10] = a[1]  & b[9];
assign y9[11] = a[2]  & b[9];
assign y9[12] = a[3]  & b[9];
assign y9[13] = a[4]  & b[9];
assign y9[14] = a[5]  & b[9];
assign y9[15] = a[6]  & b[9];
assign y9[16] = a[7]  & b[9];
assign y9[17] = a[8]  & b[9];
assign y9[18] = a[9]  & b[9];
assign y9[19] = a[10] & b[9];
assign y9[20] = a[11] & b[9];
assign y9[21] = a[12] & b[9];
assign y9[22] = a[13] & b[9];
assign y9[23] = a[14] & b[9];
assign y9[24] = a[15] & b[9];
assign y9[31:25] = 7'b0;

assign y10[9:0] = 10'b0;
assign y10[10] = a[0]  & b[10];
assign y10[11] = a[1]  & b[10];
assign y10[12] = a[2]  & b[10];
assign y10[13] = a[3]  & b[10];
assign y10[14] = a[4]  & b[10];
assign y10[15] = a[5]  & b[10];
assign y10[16] = a[6]  & b[10];
assign y10[17] = a[7]  & b[10];
assign y10[18] = a[8]  & b[10];
assign y10[19] = a[9]  & b[10];
assign y10[20] = a[10] & b[10];
assign y10[21] = a[11] & b[10];
assign y10[22] = a[12] & b[10];
assign y10[23] = a[13] & b[10];
assign y10[24] = a[14] & b[10];
assign y10[25] = a[15] & b[10];
assign y10[31:26] = 6'b0;

assign y11[10:0] = 11'b0;
assign y11[11] = a[0]  & b[11];
assign y11[12] = a[1]  & b[11];
assign y11[13] = a[2]  & b[11];
assign y11[14] = a[3]  & b[11];
assign y11[15] = a[4]  & b[11];
assign y11[16] = a[5]  & b[11];
assign y11[17] = a[6]  & b[11];
assign y11[18] = a[7]  & b[11];
assign y11[19] = a[8]  & b[11];
assign y11[20] = a[9]  & b[11];
assign y11[21] = a[10] & b[11];
assign y11[22] = a[11] & b[11];
assign y11[23] = a[12] & b[11];
assign y11[24] = a[13] & b[11];
assign y11[25] = a[14] & b[11];
assign y11[26] = a[15] & b[11];
assign y11[31:27] = 5'b0;

assign y12[11:0] = 12'b0;
assign y12[12] = a[0]  & b[12];
assign y12[13] = a[1]  & b[12];
assign y12[14] = a[2]  & b[12];
assign y12[15] = a[3]  & b[12];
assign y12[16] = a[4]  & b[12];
assign y12[17] = a[5]  & b[12];
assign y12[18] = a[6]  & b[12];
assign y12[19] = a[7]  & b[12];
assign y12[20] = a[8]  & b[12];
assign y12[21] = a[9]  & b[12];
assign y12[22] = a[10] & b[12];
assign y12[23] = a[11] & b[12];
assign y12[24] = a[12] & b[12];
assign y12[25] = a[13] & b[12];
assign y12[26] = a[14] & b[12];
assign y12[27] = a[15] & b[12];
assign y12[31:28] = 4'b0;

assign y13[12:0] = 13'b0;
assign y13[13] = a[0]  & b[13];
assign y13[14] = a[1]  & b[13];
assign y13[15] = a[2]  & b[13];
assign y13[16] = a[3]  & b[13];
assign y13[17] = a[4]  & b[13];
assign y13[18] = a[5]  & b[13];
assign y13[19] = a[6]  & b[13];
assign y13[20] = a[7]  & b[13];
assign y13[21] = a[8]  & b[13];
assign y13[22] = a[9]  & b[13];
assign y13[23] = a[10] & b[13];
assign y13[24] = a[11] & b[13];
assign y13[25] = a[12] & b[13];
assign y13[26] = a[13] & b[13];
assign y13[27] = a[14] & b[13];
assign y13[28] = a[15] & b[13];
assign y13[31:29] = 3'b0;

assign y14[13:0] = 14'b0;
assign y14[14] = a[0]  & b[14];
assign y14[15] = a[1]  & b[14];
assign y14[16] = a[2]  & b[14];
assign y14[17] = a[3]  & b[14];
assign y14[18] = a[4]  & b[14];
assign y14[19] = a[5]  & b[14];
assign y14[20] = a[6]  & b[14];
assign y14[21] = a[7]  & b[14];
assign y14[22] = a[8]  & b[14];
assign y14[23] = a[9]  & b[14];
assign y14[24] = a[10] & b[14];
assign y14[25] = a[11] & b[14];
assign y14[26] = a[12] & b[14];
assign y14[27] = a[13] & b[14];
assign y14[28] = a[14] & b[14];
assign y14[29] = a[15] & b[14];
assign y14[31:30] = 2'b0;

assign y15[14:0] = 15'b0;
assign y15[15] = a[0]  & b[15];
assign y15[16] = a[1]  & b[15];
assign y15[17] = a[2]  & b[15];
assign y15[18] = a[3]  & b[15];
assign y15[19] = a[4]  & b[15];
assign y15[20] = a[5]  & b[15];
assign y15[21] = a[6]  & b[15];
assign y15[22] = a[7]  & b[15];
assign y15[23] = a[8]  & b[15];
assign y15[24] = a[9]  & b[15];
assign y15[25] = a[10] & b[15];
assign y15[26] = a[11] & b[15];
assign y15[27] = a[12] & b[15];
assign y15[28] = a[13] & b[15];
assign y15[29] = a[14] & b[15];
assign y15[30] = a[15] & b[15];
assign y15[31] = 1'b0;


modifiedAdder_32bit add0 (.Cin(1'b0), .A(y0),  .B(y1),  .Sum(s0), .Cout(cout0));
modifiedAdder_32bit add1 (.Cin(1'b0), .A(y2),  .B(y3),  .Sum(s1), .Cout(cout1));
modifiedAdder_32bit add2 (.Cin(1'b0), .A(y4),  .B(y5),  .Sum(s2), .Cout(cout2));
modifiedAdder_32bit add3 (.Cin(1'b0), .A(y6),  .B(y7),  .Sum(s3), .Cout(cout3));
modifiedAdder_32bit add4 (.Cin(1'b0), .A(y8),  .B(y9),  .Sum(s4), .Cout(cout4));
modifiedAdder_32bit add5 (.Cin(1'b0), .A(y10), .B(y11), .Sum(s5), .Cout(cout5));
modifiedAdder_32bit add6 (.Cin(1'b0), .A(y12), .B(y13), .Sum(s6), .Cout(cout6));
modifiedAdder_32bit add7 (.Cin(1'b0), .A(y14), .B(y15), .Sum(s7), .Cout(cout7));

modifiedAdder_32bit add8  (.Cin(1'b0), .A(s0), .B(s1), .Sum(s8),  .Cout(cout8));
modifiedAdder_32bit add9  (.Cin(1'b0), .A(s2), .B(s3), .Sum(s9),  .Cout(cout9));
modifiedAdder_32bit add10 (.Cin(1'b0), .A(s4), .B(s5), .Sum(s10), .Cout(cout10));
modifiedAdder_32bit add11 (.Cin(1'b0), .A(s6), .B(s7), .Sum(s11), .Cout(cout11));

modifiedAdder_32bit add12 (.Cin(1'b0), .A(s8), .B(s9),  .Sum(s12), .Cout(cout12));
modifiedAdder_32bit add13 (.Cin(1'b0), .A(s10), .B(s11), .Sum(s13), .Cout(cout13));

modifiedAdder_32bit add14 (.Cin(1'b0), .A(s12), .B(s13), .Sum(s14), .Cout(cout14));

endmodule
